module control_reg(output reg [28:0]cwrd,
                    input [4:0]addr,
                      input clk,reset);

reg [28:0]mem[0:25];


always @(reset)
begin
mem[0]=29'd0;
mem[1]=29'b01_01_00_0000__00_001_01_0_00_00_11_00010;
mem[2]=29'b00_10_000000__01_000_00_0_00_00_11_00011;
mem[3]=29'b00_00_000010__00_010_10_0_00_00_11_00100;
mem[4]=29'b01_00_010000__01_000_01_0_00_00_01_00101;
mem[5]=29'b10_00_01_1011__00_000_01_0_00_00_01_00110; 
mem[6]=29'b01_00_000010__00_001_00_0_00_01_10_00111;
mem[7]=29'b00_11_000000__10_000_00_0_01_10_00_00000;
mem[8]=29'b01_01_000000__00_001_00_0_00_01_11_00111;
mem[9]=29'b01_01_010001__00_001_01_0_00_01_11_01010;
mem[10]=29'b00_11_100000__10_011_00_0_01_10_00_00000;
mem[11]=29'b10_00_110011__00_011_00_1_00_00_11_01000;
mem[12]=29'b01_01_010000__00_001_10_0_00_01_11_01010;
mem[13]=29'b00_00_000011__00_100_10_0_00_00_11_01110;
mem[14]=29'b10_00_110000__01_000_00_1_00_00_11_01000;
mem[15]=29'b01_01_011001__00_001_00_0_00_01_11_01010;
mem[16]=29'b01_01_010110__00_001_00_0_00_01_11_01010;
mem[17]=29'b00_00_000010__00_101_00_0_00_00_11_10010;
mem[18]=29'b10_00_000111__10_000_00_1_00_00_11_01000;
mem[19]=29'b00_00_001011__00_100_00_0_00_00_11_10100;
mem[20]=29'b01_01_000100__10_001_00_0_00_01_11_00111;
mem[21]=29'b01_00_000010__00_001_01_0_00_00_11_10110;
mem[22]=29'b00_00_001101__01_000_10_0_00_00_11_00111;
mem[23]=29'b01_01_00_0000_00_001_00_0_00_01_11_11000;
mem[24]=29'b00_10_00_0000_01_000_00_0_01_10_00_11001;
end


always @(posedge clk)
begin
    if (reset)
    begin
    cwrd=mem[5'b01000];
    end
    
    else
    if (addr <= 5'd24 && addr >= 5'd0 )
         cwrd=mem[addr];

end
endmodule
